library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use work.emp_data_types.all;

entity jet_ip_wrapper is
  port (
    clk: in std_logic;
    rst: in std_logic;
    start: in std_logic;
    input: in ldata(71 downto 0);
    done: out std_logic;
    idle: out std_logic;
    ready: out std_logic;
    output : out ldata(71 downto 0)
    );
  
end jet_ip_wrapper;

architecture rtl of jet_ip_wrapper is
  
begin

  s2pfjet_algo : entity work.hls_delay_0
    port map (
      ap_clk => clk,
      ap_rst => rst,
      ap_start => start, -- ??
      ap_done => done, -- ??
      ap_idle => idle, -- ??
      ap_ready => ready, -- ??
      inData_0 => input(0).data(7 downto 0),
      inData_1 => input(1).data(7 downto 0),
      inData_2 => input(2).data(7 downto 0),
      inData_3 => input(3).data(7 downto 0),
      inData_4 => input(4).data(7 downto 0),
      inData_5 => input(5).data(7 downto 0),
      inData_6 => input(6).data(7 downto 0),
      inData_7 => input(7).data(7 downto 0),
      inData_8 => input(8).data(7 downto 0),
      inData_9 => input(9).data(7 downto 0),
      inData_10 => input(10).data(7 downto 0),
      inData_11 => input(11).data(7 downto 0),
      inData_12 => input(12).data(7 downto 0),
      inData_13 => input(13).data(7 downto 0),
      inData_14 => input(14).data(7 downto 0),
      inData_15 => input(15).data(7 downto 0),
      inData_16 => input(16).data(7 downto 0),
      inData_17 => input(17).data(7 downto 0),
      inData_18 => input(18).data(7 downto 0),
      inData_19 => input(19).data(7 downto 0),
      inData_20 => input(20).data(7 downto 0),
      inData_21 => input(21).data(7 downto 0),
      inData_22 => input(22).data(7 downto 0),
      inData_23 => input(23).data(7 downto 0),
      inData_24 => input(24).data(7 downto 0),
      inData_25 => input(25).data(7 downto 0),
      inData_26 => input(26).data(7 downto 0),
      inData_27 => input(27).data(7 downto 0),
      inData_28 => input(28).data(7 downto 0),
      inData_29 => input(29).data(7 downto 0),
      inData_30 => input(30).data(7 downto 0),
      inData_31 => input(31).data(7 downto 0),
      inData_32 => input(32).data(7 downto 0),
      inData_33 => input(33).data(7 downto 0),
      inData_34 => input(34).data(7 downto 0),
      inData_35 => input(35).data(7 downto 0),
      inData_36 => input(36).data(7 downto 0),
      inData_37 => input(37).data(7 downto 0),
      inData_38 => input(38).data(7 downto 0),
      inData_39 => input(39).data(7 downto 0),
      inData_40 => input(40).data(7 downto 0),
      inData_41 => input(41).data(7 downto 0),
      inData_42 => input(42).data(7 downto 0),
      inData_43 => input(43).data(7 downto 0),
      inData_44 => input(44).data(7 downto 0),
      inData_45 => input(45).data(7 downto 0),
      inData_46 => input(46).data(7 downto 0),
      inData_47 => input(47).data(7 downto 0),
      inData_48 => input(48).data(7 downto 0),
      inData_49 => input(49).data(7 downto 0),
      inData_50 => input(50).data(7 downto 0),
      inData_51 => input(51).data(7 downto 0),
      inData_52 => input(52).data(7 downto 0),
      inData_53 => input(53).data(7 downto 0),
      inData_54 => input(54).data(7 downto 0),
      inData_55 => input(55).data(7 downto 0),
      inData_56 => input(56).data(7 downto 0),
      inData_57 => input(57).data(7 downto 0),
      inData_58 => input(58).data(7 downto 0),
      inData_59 => input(59).data(7 downto 0),
      inData_60 => input(60).data(7 downto 0),
      inData_61 => input(61).data(7 downto 0),
      inData_62 => input(62).data(7 downto 0),
      inData_63 => input(63).data(7 downto 0),
      inData_64 => input(64).data(7 downto 0),
      inData_65 => input(65).data(7 downto 0),
      inData_66 => input(66).data(7 downto 0),
      inData_67 => input(67).data(7 downto 0),
      inData_68 => input(68).data(7 downto 0),
      inData_69 => input(69).data(7 downto 0),
      inData_70 => input(70).data(7 downto 0),
      inData_71 => input(71).data(7 downto 0),

      outData_0 => output(0).data(7 downto 0),
      outData_1 => output(1).data(7 downto 0),
      outData_2 => output(2).data(7 downto 0),
      outData_3 => output(3).data(7 downto 0),
      outData_4 => output(4).data(7 downto 0),
      outData_5 => output(5).data(7 downto 0),
      outData_6 => output(6).data(7 downto 0),
      outData_7 => output(7).data(7 downto 0),
      outData_8 => output(8).data(7 downto 0),
      outData_9 => output(9).data(7 downto 0),
      outData_10 => output(10).data(7 downto 0),
      outData_11 => output(11).data(7 downto 0),
      outData_12 => output(12).data(7 downto 0),
      outData_13 => output(13).data(7 downto 0),
      outData_14 => output(14).data(7 downto 0),
      outData_15 => output(15).data(7 downto 0),
      outData_16 => output(16).data(7 downto 0),
      outData_17 => output(17).data(7 downto 0),
      outData_18 => output(18).data(7 downto 0),
      outData_19 => output(19).data(7 downto 0),
      outData_20 => output(20).data(7 downto 0),
      outData_21 => output(21).data(7 downto 0),
      outData_22 => output(22).data(7 downto 0),
      outData_23 => output(23).data(7 downto 0),
      outData_24 => output(24).data(7 downto 0),
      outData_25 => output(25).data(7 downto 0),
      outData_26 => output(26).data(7 downto 0),
      outData_27 => output(27).data(7 downto 0),
      outData_28 => output(28).data(7 downto 0),
      outData_29 => output(29).data(7 downto 0),
      outData_30 => output(30).data(7 downto 0),
      outData_31 => output(31).data(7 downto 0),
      outData_32 => output(32).data(7 downto 0),
      outData_33 => output(33).data(7 downto 0),
      outData_34 => output(34).data(7 downto 0),
      outData_35 => output(35).data(7 downto 0),
      outData_36 => output(36).data(7 downto 0),
      outData_37 => output(37).data(7 downto 0),
      outData_38 => output(38).data(7 downto 0),
      outData_39 => output(39).data(7 downto 0),
      outData_40 => output(40).data(7 downto 0),
      outData_41 => output(41).data(7 downto 0),
      outData_42 => output(42).data(7 downto 0),
      outData_43 => output(43).data(7 downto 0),
      outData_44 => output(44).data(7 downto 0),
      outData_45 => output(45).data(7 downto 0),
      outData_46 => output(46).data(7 downto 0),
      outData_47 => output(47).data(7 downto 0),
      outData_48 => output(48).data(7 downto 0),
      outData_49 => output(49).data(7 downto 0),
      outData_50 => output(50).data(7 downto 0),
      outData_51 => output(51).data(7 downto 0),
      outData_52 => output(52).data(7 downto 0),
      outData_53 => output(53).data(7 downto 0),
      outData_54 => output(54).data(7 downto 0),
      outData_55 => output(55).data(7 downto 0),
      outData_56 => output(56).data(7 downto 0),
      outData_57 => output(57).data(7 downto 0),
      outData_58 => output(58).data(7 downto 0),
      outData_59 => output(59).data(7 downto 0),
      outData_60 => output(60).data(7 downto 0),
      outData_61 => output(61).data(7 downto 0),
      outData_62 => output(62).data(7 downto 0),
      outData_63 => output(63).data(7 downto 0),
      outData_64 => output(64).data(7 downto 0),
      outData_65 => output(65).data(7 downto 0),
      outData_66 => output(66).data(7 downto 0),
      outData_67 => output(67).data(7 downto 0),
      outData_68 => output(68).data(7 downto 0),
      outData_69 => output(69).data(7 downto 0),
      outData_70 => output(70).data(7 downto 0),
      outData_71 => output(71).data(7 downto 0)
      );

end rtl;

