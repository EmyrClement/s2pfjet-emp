library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use work.emp_data_types.all;

entity jet_ip_wrapper is
  port (
    clk: in std_logic;
    rst: in std_logic;
    start: in std_logic;
    input: in ldata(71 downto 0);
    done: out std_logic;
    idle: out std_logic;
    ready: out std_logic;
    output : out ldata(71 downto 0)
    );
  
end jet_ip_wrapper;

architecture rtl of jet_ip_wrapper is
  
begin

  s2pfjet_algo : entity work.hls_delay_0
    port map (
      ap_clk => clk,
      ap_rst => rst,
      ap_start => start, -- ??
      ap_done => done, -- ??
      ap_idle => idle, -- ??
      ap_ready => ready, -- ??
      inData_0_V => input(0).data,
      inData_1_V => input(1).data,
      inData_2_V => input(2).data,
      inData_3_V => input(3).data,
      inData_4_V => input(4).data,
      inData_5_V => input(5).data,
      inData_6_V => input(6).data,
      inData_7_V => input(7).data,
      inData_8_V => input(8).data,
      inData_9_V => input(9).data,
      inData_10_V => input(10).data,
      inData_11_V => input(11).data,
      inData_12_V => input(12).data,
      inData_13_V => input(13).data,
      inData_14_V => input(14).data,
      inData_15_V => input(15).data,
      inData_16_V => input(16).data,
      inData_17_V => input(17).data,
      inData_18_V => input(18).data,
      inData_19_V => input(19).data,
      inData_20_V => input(20).data,
      inData_21_V => input(21).data,
      inData_22_V => input(22).data,
      inData_23_V => input(23).data,
      inData_24_V => input(24).data,
      inData_25_V => input(25).data,
      inData_26_V => input(26).data,
      inData_27_V => input(27).data,
      inData_28_V => input(28).data,
      inData_29_V => input(29).data,
      inData_30_V => input(30).data,
      inData_31_V => input(31).data,
      inData_32_V => input(32).data,
      inData_33_V => input(33).data,
      inData_34_V => input(34).data,
      inData_35_V => input(35).data,
      inData_36_V => input(36).data,
      inData_37_V => input(37).data,
      inData_38_V => input(38).data,
      inData_39_V => input(39).data,
      inData_40_V => input(40).data,
      inData_41_V => input(41).data,
      inData_42_V => input(42).data,
      inData_43_V => input(43).data,
      inData_44_V => input(44).data,
      inData_45_V => input(45).data,
      inData_46_V => input(46).data,
      inData_47_V => input(47).data,
      inData_48_V => input(48).data,
      inData_49_V => input(49).data,
      inData_50_V => input(50).data,
      inData_51_V => input(51).data,
      inData_52_V => input(52).data,
      inData_53_V => input(53).data,
      inData_54_V => input(54).data,
      inData_55_V => input(55).data,
      inData_56_V => input(56).data,
      inData_57_V => input(57).data,
      inData_58_V => input(58).data,
      inData_59_V => input(59).data,
      inData_60_V => input(60).data,
      inData_61_V => input(61).data,
      inData_62_V => input(62).data,
      inData_63_V => input(63).data,
      inData_64_V => input(64).data,
      inData_65_V => input(65).data,
      inData_66_V => input(66).data,
      inData_67_V => input(67).data,
      inData_68_V => input(68).data,
      inData_69_V => input(69).data,
      inData_70_V => input(70).data,
      inData_71_V => input(71).data,

      outData_0_V => output(0).data,
      outData_1_V => output(1).data,
      outData_2_V => output(2).data,
      outData_3_V => output(3).data,
      outData_4_V => output(4).data,
      outData_5_V => output(5).data,
      outData_6_V => output(6).data,
      outData_7_V => output(7).data,
      outData_8_V => output(8).data,
      outData_9_V => output(9).data,
      outData_10_V => output(10).data,
      outData_11_V => output(11).data,
      outData_12_V => output(12).data,
      outData_13_V => output(13).data,
      outData_14_V => output(14).data,
      outData_15_V => output(15).data,
      outData_16_V => output(16).data,
      outData_17_V => output(17).data,
      outData_18_V => output(18).data,
      outData_19_V => output(19).data,
      outData_20_V => output(20).data,
      outData_21_V => output(21).data,
      outData_22_V => output(22).data,
      outData_23_V => output(23).data,
      outData_24_V => output(24).data,
      outData_25_V => output(25).data,
      outData_26_V => output(26).data,
      outData_27_V => output(27).data,
      outData_28_V => output(28).data,
      outData_29_V => output(29).data,
      outData_30_V => output(30).data,
      outData_31_V => output(31).data,
      outData_32_V => output(32).data,
      outData_33_V => output(33).data,
      outData_34_V => output(34).data,
      outData_35_V => output(35).data,
      outData_36_V => output(36).data,
      outData_37_V => output(37).data,
      outData_38_V => output(38).data,
      outData_39_V => output(39).data,
      outData_40_V => output(40).data,
      outData_41_V => output(41).data,
      outData_42_V => output(42).data,
      outData_43_V => output(43).data,
      outData_44_V => output(44).data,
      outData_45_V => output(45).data,
      outData_46_V => output(46).data,
      outData_47_V => output(47).data,
      outData_48_V => output(48).data,
      outData_49_V => output(49).data,
      outData_50_V => output(50).data,
      outData_51_V => output(51).data,
      outData_52_V => output(52).data,
      outData_53_V => output(53).data,
      outData_54_V => output(54).data,
      outData_55_V => output(55).data,
      outData_56_V => output(56).data,
      outData_57_V => output(57).data,
      outData_58_V => output(58).data,
      outData_59_V => output(59).data,
      outData_60_V => output(60).data,
      outData_61_V => output(61).data,
      outData_62_V => output(62).data,
      outData_63_V => output(63).data,
      outData_64_V => output(64).data,
      outData_65_V => output(65).data,
      outData_66_V => output(66).data,
      outData_67_V => output(67).data,
      outData_68_V => output(68).data,
      outData_69_V => output(69).data,
      outData_70_V => output(70).data,
      outData_71_V => output(71).data
      );

end rtl;

